module vopengl

#flag -Ivendor/include

