module main
#flag -Ivendor/include
#flag -Lvendor/lib/libglfw3.a
#include "glad/glad.h"
#include "GLFW/glfw3.h"


fn main() {
	println('Hello World!')
}
