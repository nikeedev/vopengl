module vopengl

[typedef]
pub type GLhandleARB = &voidptr
