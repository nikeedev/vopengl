module main
import vopengl


fn run() {
	vopengl.
}
