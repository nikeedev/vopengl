module vopengl

[typedef]
pub type GLhandleARB = u32
